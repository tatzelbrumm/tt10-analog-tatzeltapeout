MACRO tatzeltapeout_tile
  CLASS BLOCK ;
  FOREIGN tatzeltapeout_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 225.760 ;
  OBS
      LAYER met4 ;
        RECT 58.000 1.000 138.560 1.500 ;
  END
END tatzeltapeout_tile
END LIBRARY

