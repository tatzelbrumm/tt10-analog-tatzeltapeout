MACRO tatzeltapeout_tile
  CLASS BLOCK ;
  FOREIGN tatzeltapeout_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  OBS
      LAYER met4 ;
        RECT 73.530 1.000 153.710 1.500 ;
  END
END tatzeltapeout_tile
END LIBRARY

