magic
tech sky130A
timestamp 1740695003
<< metal4 >>
rect 13239 100 15281 150
<< properties >>
string FIXED_BBOX 0 0 33488 22576
<< end >>
