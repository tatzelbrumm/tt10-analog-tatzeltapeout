magic
tech sky130A
timestamp 1740695003
<< isosubstrate >>
rect 0 0 14536 22576
<< metal4 >>
rect 5800 100 13856 150
<< properties >>
string FIXED_BBOX 0 0 14536 22576
<< end >>
